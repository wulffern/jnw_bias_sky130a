magic
tech sky130A
magscale 1 2
timestamp 1755986400
<< checkpaint >>
rect 0 0 28354 10560
<< m3 >>
rect 8552 4874 12352 5074
rect 8992 4434 9192 9594
rect 10352 4434 10552 9594
rect 11712 4434 11912 9594
rect 8552 6234 12352 6434
rect 8992 4434 9192 9594
rect 10352 4434 10552 9594
rect 11712 4434 11912 9594
rect 8552 7594 12352 7794
rect 8992 4434 9192 9594
rect 10352 4434 10552 9594
rect 11712 4434 11912 9594
rect 8552 8954 9632 9154
rect 8992 4434 9192 9594
<< m4 >>
rect 8552 4874 12352 5074
rect 8992 4434 9192 9594
rect 10352 4434 10552 9594
rect 11712 4434 11912 9594
rect 8552 6234 12352 6434
rect 8992 4434 9192 9594
rect 10352 4434 10552 9594
rect 11712 4434 11912 9594
rect 8552 7594 12352 7794
rect 8992 4434 9192 9594
rect 10352 4434 10552 9594
rect 11712 4434 11912 9594
rect 8552 8954 9632 9154
rect 8992 4434 9192 9594
use JNWBIAS_OTACM xaota6 ../JNW_BIAS_SKY130A
transform 1 0 0 0 1 0
box 0 0 6800 10000
use JNWATR_PCH_4CTAPBOT xb1<0>_BOT ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 0
box 7100 0 8252 480
use JNWATR_PCH_4C5F0 xb1<0> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 480
box 7100 480 8252 1280
use JNWATR_PCH_4C5F0 xb1<1> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 1280
box 7100 1280 8252 2080
use JNWATR_PCH_4C5F0 xb1<2> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 2080
box 7100 2080 8252 2880
use JNWATR_PCH_4C5F0 xb1<3> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 2880
box 7100 2880 8252 3680
use JNWATR_PCH_4C5F0 xb3<0> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 3680
box 7100 3680 8252 4480
use JNWATR_PCH_4C5F0 xb3<1> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 4480
box 7100 4480 8252 5280
use JNWATR_PCH_4C5F0 xb3<2> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 5280
box 7100 5280 8252 6080
use JNWATR_PCH_4C5F0 xb3<3> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 6080
box 7100 6080 8252 6880
use JNWATR_PCH_4C5F0 xb7<0> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 6880
box 7100 6880 8252 7680
use JNWATR_PCH_4C5F0 xb7<1> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 7680
box 7100 7680 8252 8480
use JNWATR_PCH_4C5F0 xb7<2> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 8480
box 7100 8480 8252 9280
use JNWATR_PCH_4C5F0 xb7<3> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 9280
box 7100 9280 8252 10080
use JNWATR_PCH_4CTAPTOP xb7<3>_TOP ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 10080
box 7100 10080 8252 10560
use JNWBIAS_BIPOLAR xbc1 ../JNW_BIAS_SKY130A
transform 1 0 8552 0 1 0
box 8552 0 12986 4434
use JNWTR_CAPX1 xbc2<0> ../JNW_TR_SKY130A
transform 1 0 8552 0 1 4434
box 8552 4434 9632 5514
use JNWTR_CAPX1 xbc2<1> ../JNW_TR_SKY130A
transform 1 0 9912 0 1 4434
box 9912 4434 10992 5514
use JNWTR_CAPX1 xbc2<2> ../JNW_TR_SKY130A
transform 1 0 11272 0 1 4434
box 11272 4434 12352 5514
use JNWTR_CAPX1 xbc2<3> ../JNW_TR_SKY130A
transform 1 0 8552 0 1 5794
box 8552 5794 9632 6874
use JNWTR_CAPX1 xbc2<4> ../JNW_TR_SKY130A
transform 1 0 9912 0 1 5794
box 9912 5794 10992 6874
use JNWTR_CAPX1 xbc2<5> ../JNW_TR_SKY130A
transform 1 0 11272 0 1 5794
box 11272 5794 12352 6874
use JNWTR_CAPX1 xbc2<6> ../JNW_TR_SKY130A
transform 1 0 8552 0 1 7154
box 8552 7154 9632 8234
use JNWTR_CAPX1 xbc2<7> ../JNW_TR_SKY130A
transform 1 0 9912 0 1 7154
box 9912 7154 10992 8234
use JNWTR_CAPX1 xbc2<8> ../JNW_TR_SKY130A
transform 1 0 11272 0 1 7154
box 11272 7154 12352 8234
use JNWTR_CAPX1 xbc2<9> ../JNW_TR_SKY130A
transform 1 0 8552 0 1 8514
box 8552 8514 9632 9594
use JNWTR_RPPO8 xc11 ../JNW_TR_SKY130A
transform 1 0 13186 0 1 0
box 13186 0 15930 3440
use JNWTR_RPPO16 xc12 ../JNW_TR_SKY130A
transform 1 0 13186 0 1 3440
box 13186 3440 17658 6880
use JNWTR_RPPO16 xc9 ../JNW_TR_SKY130A
transform 1 0 13186 0 1 6880
box 13186 6880 17658 10320
use JNWTR_RPPO8 xd10 ../JNW_TR_SKY130A
transform 1 0 17858 0 1 0
box 17858 0 20602 3440
use JNWTR_RPPO16 xd13 ../JNW_TR_SKY130A
transform 1 0 17858 0 1 3440
box 17858 3440 22330 6880
use JNWTR_RPPO16 xd7 ../JNW_TR_SKY130A
transform 1 0 17858 0 1 6880
box 17858 6880 22330 10320
use JNWTR_RPPO4 xe2 ../JNW_TR_SKY130A
transform 1 0 22530 0 1 0
box 22530 0 24410 3440
use JNWTR_RPPO16 xe3 ../JNW_TR_SKY130A
transform 1 0 22530 0 1 3440
box 22530 3440 27002 6880
use JNWTR_RPPO2 xe8 ../JNW_TR_SKY130A
transform 1 0 22530 0 1 6880
box 22530 6880 23978 10320
use JNWATR_NCH_4CTAPBOT xf4_BOT ../JNW_ATR_SKY130A
transform 1 0 27202 0 1 0
box 27202 0 28354 480
use JNWATR_NCH_4C5F0 xf4 ../JNW_ATR_SKY130A
transform 1 0 27202 0 1 480
box 27202 480 28354 1280
use JNWATR_NCH_4CTAPTOP xf4_TOP ../JNW_ATR_SKY130A
transform 1 0 27202 0 1 1280
box 27202 1280 28354 1760
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 28354 10560
<< end >>
