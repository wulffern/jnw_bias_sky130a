magic
tech sky130A
magscale 1 2
timestamp 1756047484
<< locali >>
rect -400 4000 -120 5240
rect 900 4000 1720 6840
rect -400 3600 1720 4000
rect -400 3200 10700 3600
rect -400 0 -120 3200
rect 1160 3100 10700 3200
rect 100 2960 500 3000
rect 100 2720 180 2960
rect 420 2720 500 2960
rect 100 2700 500 2720
rect 1160 0 1500 3100
rect 3180 0 3480 3100
rect 6060 0 6340 3100
rect -400 -400 11600 0
<< viali >>
rect 1980 6320 2220 6560
rect 5486 6326 5714 6554
rect 6580 6320 6820 6560
rect 10074 6386 10302 6614
rect 180 2720 420 2960
rect 596 2720 836 2960
rect 1786 2726 2014 2954
rect 2676 2720 2916 2960
rect 3786 2726 4014 2954
rect 5540 2720 5780 2960
rect 6586 2726 6814 2954
rect 10068 2720 10308 2960
<< metal1 >>
rect 1974 7580 1980 7820
rect 2220 7580 2226 7820
rect 1980 6600 2220 7580
rect 10000 6614 10400 6700
rect 1900 6560 2300 6600
rect 1900 6320 1980 6560
rect 2220 6320 2300 6560
rect 1900 6300 2300 6320
rect 5400 6560 5800 6600
rect 6500 6560 6900 6600
rect 5400 6554 6580 6560
rect 5400 6326 5486 6554
rect 5714 6326 6580 6554
rect 5400 6320 6580 6326
rect 6820 6320 6900 6560
rect 5400 6300 5800 6320
rect 6500 6300 6900 6320
rect 10000 6386 10074 6614
rect 10302 6386 10400 6614
rect 10000 6300 10400 6386
rect 180 3000 420 4720
rect 10068 3100 10308 6300
rect 100 2960 500 3000
rect 100 2720 180 2960
rect 420 2720 500 2960
rect 100 2700 500 2720
rect 580 2960 1000 3100
rect 1700 2960 2100 3100
rect 580 2720 596 2960
rect 836 2954 2100 2960
rect 836 2726 1786 2954
rect 2014 2726 2100 2954
rect 836 2720 2100 2726
rect 580 2700 1000 2720
rect 1700 2700 2100 2720
rect 2600 2960 3000 3000
rect 3700 2960 4100 3000
rect 2600 2720 2676 2960
rect 2916 2954 4100 2960
rect 2916 2726 3786 2954
rect 4014 2726 4100 2954
rect 2916 2720 4100 2726
rect 2600 2600 3000 2720
rect 3700 2600 4100 2720
rect 5500 2960 5900 3100
rect 6500 2960 6900 3100
rect 5500 2720 5540 2960
rect 5780 2954 6900 2960
rect 5780 2726 6586 2954
rect 6814 2726 6900 2954
rect 5780 2720 6900 2726
rect 5500 2700 5900 2720
rect 6500 2700 6900 2720
rect 10000 2960 10400 3100
rect 10000 2720 10068 2960
rect 10308 2720 10400 2960
rect 10000 2700 10400 2720
<< via1 >>
rect 1980 7580 2220 7820
<< metal2 >>
rect 1980 7823 2220 7826
rect -322 7820 2223 7823
rect -322 7580 1980 7820
rect 2220 7580 2223 7820
rect -322 7578 2223 7580
rect 1980 7574 2220 7578
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1734020192
transform 1 0 -200 0 1 3800
box 0 0 1340 1340
use JNWTR_RPPO2  xa1 ../JNW_TR_SKY130A
timestamp 1755255778
transform 1 0 -200 0 1 -200
box 0 0 1448 3440
use JNWTR_RPPO4  xb1 ../JNW_TR_SKY130A
timestamp 1755333658
transform 1 0 1400 0 1 -200
box 0 0 1880 3440
use JNWTR_RPPO8  xc1 ../JNW_TR_SKY130A
timestamp 1755344196
transform 1 0 3400 0 1 -200
box 0 0 2744 3440
use JNWTR_RPPO16  xd3_0 ../JNW_TR_SKY130A
timestamp 1756043915
transform -1 0 6072 0 1 3400
box 0 0 4472 3440
use JNWTR_RPPO16  xd3_1
timestamp 1756043915
transform -1 0 10672 0 1 3400
box 0 0 4472 3440
use JNWTR_RPPO16  xd3_2
timestamp 1756043915
transform 1 0 6200 0 1 -200
box 0 0 4472 3440
<< labels >>
flabel locali -400 -400 11600 0 0 FreeSans 1600 0 0 0 VSS
port 0 nsew
flabel metal2 -322 7578 1980 7823 0 FreeSans 1600 0 0 0 VREF
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 6472 3440
<< end >>
