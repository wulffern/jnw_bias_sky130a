magic
tech sky130A
magscale 1 2
timestamp 1755335025
<< psubdiff >>
rect -117 4283 -57 4317
rect 4257 4283 4317 4317
rect -117 4257 -83 4283
rect -117 -83 -83 -57
rect 4283 4257 4317 4283
rect 4283 -83 4317 -57
rect -117 -117 -57 -83
rect 4257 -117 4317 -83
<< psubdiffcont >>
rect -57 4283 4257 4317
rect -117 -57 -83 4257
rect 4283 -57 4317 4257
rect -57 -117 4257 -83
<< locali >>
rect -117 4283 -57 4317
rect 4257 4283 4317 4317
rect -117 4257 -83 4283
rect 4283 4257 4317 4283
rect -117 -83 -83 -57
rect 20 3940 4160 4160
rect 20 3080 240 3940
rect 1100 3080 1660 3940
rect 2520 3080 3080 3940
rect 3940 3080 4160 3940
rect 20 2520 4160 3080
rect 20 1660 240 2520
rect 1100 1660 1660 2520
rect 2520 1660 3080 2520
rect 3940 1660 4160 2520
rect 20 1100 4160 1660
rect 20 240 240 1100
rect 1100 240 1660 1100
rect 2520 240 3080 1100
rect 3940 240 4160 1100
rect 20 -83 4160 240
rect 4283 -83 4317 -57
rect -117 -117 -57 -83
rect 4257 -117 4317 -83
<< metal1 >>
rect 300 3100 3900 3900
rect 300 1000 1100 3100
rect 1700 1700 2500 2500
rect 3100 1000 3900 3100
rect 300 300 3900 1000
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 2 1420 0 2 1420
timestamp 1755333750
transform 1 0 0 0 1 0
box 0 0 1340 1340
<< labels >>
flabel metal1 1700 1700 2500 2500 0 FreeSans 1600 0 0 0 VD1
port 0 nsew
flabel metal1 300 3100 3900 3900 0 FreeSans 1600 0 0 0 VD2
port 1 nsew
flabel locali s 20 -100 4160 140 0 FreeSans 1600 0 0 0 VSS
port 2 nsew
<< end >>
