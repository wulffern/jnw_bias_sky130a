magic
tech sky130A
magscale 1 2
timestamp 1755460977
<< locali >>
rect 3908 10000 4290 10002
rect 0 9921 9600 10000
rect 0 9890 2982 9921
rect 0 9710 678 9890
rect 858 9886 2982 9890
rect 858 9885 2854 9886
rect 858 9710 1830 9885
rect 0 9705 1830 9710
rect 2010 9834 2854 9885
rect 2906 9834 2982 9886
rect 2010 9741 2982 9834
rect 3162 9908 9600 9921
rect 3162 9902 9608 9908
rect 3162 9898 8298 9902
rect 3162 9741 3366 9898
rect 2010 9718 3366 9741
rect 3546 9718 8298 9898
rect 2010 9705 8298 9718
rect 0 9698 8298 9705
rect 8502 9698 9608 9902
rect 0 9692 9608 9698
rect 0 9600 9600 9692
rect 0 9592 400 9600
rect 0 9492 1500 9592
rect 3162 9580 3936 9600
rect 0 4300 400 9492
rect 14800 6200 15200 10000
rect 0 400 400 3800
rect 580 2700 820 2780
rect 580 1100 840 1180
rect 3600 400 3900 3500
rect 5020 3460 5340 3480
rect 5020 3220 5040 3460
rect 5280 3220 5340 3460
rect 5020 3200 5340 3220
rect 5600 400 5900 4700
rect 14800 400 15200 6000
rect 0 294 15200 400
rect 0 66 3046 294
rect 3274 66 15200 294
rect 0 0 15200 66
<< viali >>
rect 678 9710 858 9890
rect 1830 9705 2010 9885
rect 2854 9834 2906 9886
rect 2982 9741 3162 9921
rect 3366 9718 3546 9898
rect 8298 9698 8502 9902
rect 2170 3250 2350 3430
rect 3040 3220 3280 3460
rect 4190 3270 4370 3450
rect 5040 3220 5280 3460
rect 6146 3226 6374 3454
rect 7970 3250 8150 3430
rect 3046 66 3274 294
<< metal1 >>
rect 2976 9921 3168 9933
rect 672 9890 864 9902
rect 672 9710 678 9890
rect 858 9710 864 9890
rect 544 9532 608 9538
rect 608 9468 614 9524
rect 544 9460 614 9468
rect 544 4332 608 9460
rect 672 4904 864 9710
rect 1824 9885 2016 9897
rect 1824 9705 1830 9885
rect 2010 9705 2016 9885
rect 2842 9886 2918 9892
rect 2842 9834 2854 9886
rect 2906 9834 2918 9886
rect 2842 9828 2918 9834
rect 1050 8676 1056 8868
rect 1248 8676 1254 8868
rect 1050 7796 1056 7988
rect 1248 7796 1254 7988
rect 1040 7524 1260 7532
rect 1040 7332 1056 7524
rect 1248 7332 1260 7524
rect 1040 7312 1260 7332
rect 1056 6816 1248 6822
rect 1056 6224 1248 6624
rect 1696 4782 1760 8683
rect 1824 4889 2016 9705
rect 2208 6822 2400 8839
rect 2193 6816 2400 6822
rect 2385 6624 2400 6816
rect 2193 6618 2400 6624
rect 2208 4949 2400 6618
rect 2848 5971 2912 9828
rect 2976 9741 2982 9921
rect 3162 9741 3168 9921
rect 2976 4717 3168 9741
rect 3360 9898 3552 9910
rect 3360 9718 3366 9898
rect 3546 9718 3552 9898
rect 3360 5791 3552 9718
rect 7992 9908 8208 9914
rect 8208 9902 8514 9908
rect 8208 9698 8298 9902
rect 8502 9698 8514 9902
rect 8208 9692 8514 9698
rect 7992 9686 8208 9692
rect 14352 9596 14544 9602
rect 14352 9020 14544 9404
rect 14352 7844 14544 8760
rect 3960 7524 4200 7540
rect 3960 7332 3985 7524
rect 4177 7332 4200 7524
rect 3960 7320 4200 7332
rect 3648 6818 3840 6824
rect 3648 5188 3840 6626
rect 3360 4996 3840 5188
rect 544 4262 608 4268
rect 1468 4332 1532 4338
rect 1468 4262 1532 4268
rect 1696 4312 1760 4616
rect 2848 4312 2912 4671
rect 1696 4262 2912 4312
rect 1468 4248 2912 4262
rect 1468 4198 1760 4248
rect 1056 4116 1248 4122
rect 672 3776 864 3782
rect 672 2724 864 3584
rect 1056 2772 1248 3924
rect 1468 2232 1532 4198
rect 3985 4115 4177 7320
rect 5998 6904 6004 7096
rect 6196 6904 6202 7096
rect 8644 6816 8836 6822
rect 8836 6624 8996 6816
rect 8644 6618 8836 6624
rect 3985 3917 4177 3923
rect 4184 3776 4376 3782
rect 3020 3460 3340 3480
rect 1168 2168 1532 2232
rect 2164 3430 2356 3442
rect 2164 3250 2170 3430
rect 2350 3250 2356 3430
rect 540 1580 604 2064
rect 678 1624 684 1816
rect 876 1624 882 1816
rect 1040 1500 1260 1520
rect 1040 1308 1056 1500
rect 1248 1308 1260 1500
rect 1040 1300 1260 1308
rect 672 1116 864 1122
rect 672 918 864 924
rect 2164 1116 2356 3250
rect 3020 3220 3040 3460
rect 3280 3220 3340 3460
rect 4184 3450 4376 3584
rect 6104 3776 6296 5596
rect 10304 4116 10496 4122
rect 7958 3924 7964 4116
rect 8156 3924 8162 4116
rect 10496 3924 10656 4116
rect 6104 3578 6296 3584
rect 4184 3270 4190 3450
rect 4370 3270 4376 3450
rect 4184 3258 4376 3270
rect 5020 3460 5340 3480
rect 6140 3460 6460 3480
rect 5020 3220 5040 3460
rect 5280 3454 6460 3460
rect 5280 3226 6146 3454
rect 6374 3226 6460 3454
rect 7964 3430 8156 3924
rect 10304 3918 10496 3924
rect 7964 3250 7970 3430
rect 8150 3250 8156 3430
rect 7964 3238 8156 3250
rect 5280 3220 6460 3226
rect 3034 3214 3286 3220
rect 2164 918 2356 924
rect 3040 294 3280 3214
rect 5020 3200 5340 3220
rect 6140 3200 6460 3220
rect 3040 66 3046 294
rect 3274 66 3280 294
rect 3040 54 3280 66
<< via1 >>
rect 544 9468 608 9532
rect 1056 8676 1248 8868
rect 1056 7796 1248 7988
rect 1056 7332 1248 7524
rect 1056 6624 1248 6816
rect 1056 5396 1248 5588
rect 1056 4596 1248 4788
rect 2193 6624 2385 6816
rect 7992 9692 8208 9908
rect 14352 9404 14544 9596
rect 3985 7332 4177 7524
rect 3648 6626 3840 6818
rect 544 4268 608 4332
rect 1468 4268 1532 4332
rect 1056 3924 1248 4116
rect 672 3584 864 3776
rect 6004 6904 6196 7096
rect 8644 6624 8836 6816
rect 3985 3923 4177 4115
rect 4184 3584 4376 3776
rect 684 1624 876 1816
rect 1056 1308 1248 1500
rect 672 924 864 1116
rect 7964 3924 8156 4116
rect 10304 3924 10496 4116
rect 6104 3584 6296 3776
rect 2164 924 2356 1116
<< metal2 >>
rect 8697 9908 8903 9912
rect 7986 9692 7992 9908
rect 8208 9903 8908 9908
rect 8208 9697 8697 9903
rect 8903 9697 8908 9903
rect 8208 9692 8908 9697
rect 8697 9688 8903 9692
rect 6796 9600 6805 9675
rect 460 9532 6805 9600
rect 460 9524 544 9532
rect 461 9468 544 9524
rect 608 9468 6805 9532
rect 461 9460 6805 9468
rect 460 9400 6805 9460
rect 6796 9285 6805 9400
rect 7195 9600 7204 9675
rect 7195 9596 14600 9600
rect 7195 9404 14352 9596
rect 14544 9404 14600 9596
rect 7195 9400 14600 9404
rect 7195 9285 7204 9400
rect 1056 8868 1248 8874
rect 0 8676 1056 8868
rect 1056 8670 1248 8676
rect 4 7988 100 7996
rect 1056 7992 1248 7994
rect 1040 7988 1260 7992
rect 4 7804 1056 7988
rect 100 7796 1056 7804
rect 1248 7796 1260 7988
rect 1040 7772 1260 7796
rect 1040 7524 1260 7532
rect 1040 7332 1056 7524
rect 1248 7332 3985 7524
rect 4177 7332 4510 7524
rect 1040 7312 1260 7332
rect 6004 7096 6196 7102
rect 3642 6816 3648 6818
rect 1050 6624 1056 6816
rect 1248 6624 2193 6816
rect 2385 6626 3648 6816
rect 3840 6816 3846 6818
rect 6004 6816 6196 6904
rect 3840 6626 8644 6816
rect 2385 6624 8644 6626
rect 8836 6624 8842 6816
rect 4 5588 100 5596
rect 1060 5588 1280 5612
rect 4 5404 1056 5588
rect 100 5396 1056 5404
rect 1248 5396 1280 5588
rect 1060 5392 1280 5396
rect 4 4788 100 4796
rect 1040 4788 1260 4792
rect 4 4604 1056 4788
rect 100 4596 1056 4604
rect 1248 4596 1260 4788
rect 1040 4572 1260 4596
rect 538 4268 544 4332
rect 608 4268 1468 4332
rect 1532 4268 1538 4332
rect 7964 4116 8156 4122
rect 1050 3924 1056 4116
rect 1248 4115 7964 4116
rect 1248 3924 3985 4115
rect 3979 3923 3985 3924
rect 4177 3924 7964 4115
rect 8156 3924 10304 4116
rect 10496 3924 10502 4116
rect 4177 3923 4183 3924
rect 7964 3918 8156 3924
rect 666 3584 672 3776
rect 864 3584 4184 3776
rect 4376 3584 6104 3776
rect 6296 3584 7110 3776
rect 684 1816 876 1822
rect 684 1500 876 1624
rect 1040 1500 1260 1520
rect 684 1308 1056 1500
rect 1248 1308 1260 1500
rect 1040 1300 1260 1308
rect 666 924 672 1116
rect 864 924 2164 1116
rect 2356 924 2362 1116
<< via2 >>
rect 8697 9697 8903 9903
rect 6805 9285 7195 9675
<< metal3 >>
rect 8292 9907 8908 9908
rect 8287 9693 8293 9907
rect 8507 9903 8908 9907
rect 8507 9697 8697 9903
rect 8903 9697 8908 9903
rect 8507 9693 8908 9697
rect 8292 9692 8908 9693
rect 6800 9675 7200 9680
rect 6800 9285 6805 9675
rect 7195 9285 7200 9675
rect 6800 8800 7200 9285
rect 6800 8400 8000 8800
rect 6800 3800 7200 8400
rect 8200 3800 8600 9080
<< via3 >>
rect 8293 9693 8507 9907
<< metal4 >>
rect 8292 9907 8508 9908
rect 8292 9693 8293 9907
rect 8507 9693 8508 9907
rect 6800 8800 7200 9100
rect 8292 9080 8508 9693
rect 6800 8400 8000 8800
rect 6800 4000 7200 8400
rect 8200 3800 8600 9080
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 384 0 1 1540
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1740610800
transform 1 0 384 0 1 2340
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 1536 0 1 4500
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_1
timestamp 1740610800
transform 1 0 1536 0 1 5300
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_2
timestamp 1740610800
transform 1 0 1536 0 1 6100
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_3
timestamp 1740610800
transform 1 0 1536 0 1 7700
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_4
timestamp 1740610800
transform 1 0 1536 0 1 6900
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_5
timestamp 1740610800
transform 1 0 1536 0 1 8500
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_6
timestamp 1740610800
transform 1 0 2688 0 1 6100
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_7
timestamp 1740610800
transform 1 0 2688 0 1 6900
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_8
timestamp 1740610800
transform 1 0 2688 0 1 7700
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_9
timestamp 1740610800
transform 1 0 2688 0 1 8500
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_10
timestamp 1740610800
transform 1 0 2688 0 1 5300
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_11
timestamp 1740610800
transform 1 0 2688 0 1 4500
box -184 -128 1336 928
use JNWATR_PCH_4CTAPBOT  JNWATR_PCH_4CTAPBOT_0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform -1 0 2688 0 1 4039
box -184 -128 1336 608
use JNWATR_PCH_4CTAPBOT  JNWATR_PCH_4CTAPBOT_1
timestamp 1740610800
transform -1 0 3840 0 1 4039
box -184 -128 1336 608
use JNWATR_PCH_4CTAPTOP  JNWATR_PCH_4CTAPTOP_0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 1536 0 1 9300
box -184 -128 1336 608
use JNWATR_PCH_4CTAPTOP  JNWATR_PCH_4CTAPTOP_1
timestamp 1740610800
transform 1 0 2688 0 1 9300
box -184 -128 1336 608
use JNWTR_CAPX1  JNWTR_CAPX1_0 ../JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 7900 0 1 5200
box 0 0 1080 1080
use JNWTR_CAPX1  JNWTR_CAPX1_1
timestamp 1737500400
transform 1 0 6500 0 1 6600
box 0 0 1080 1080
use JNWTR_CAPX1  JNWTR_CAPX1_2
timestamp 1737500400
transform 1 0 7900 0 1 6600
box 0 0 1080 1080
use JNWTR_CAPX1  JNWTR_CAPX1_3
timestamp 1737500400
transform 1 0 6500 0 1 8000
box 0 0 1080 1080
use JNWTR_CAPX1  JNWTR_CAPX1_4
timestamp 1737500400
transform 1 0 7900 0 1 8000
box 0 0 1080 1080
use JNWTR_CAPX1  JNWTR_CAPX1_5
timestamp 1737500400
transform 1 0 7900 0 1 3800
box 0 0 1080 1080
use JNWTR_CAPX1  JNWTR_CAPX1_6
timestamp 1737500400
transform 1 0 6500 0 1 3800
box 0 0 1080 1080
use JNWTR_RPPO8  xab3 ../JNW_TR_SKY130A
timestamp 1755344196
transform 1 0 5800 0 1 300
box 0 0 2744 3440
use JNWTR_RPPO4  xac2 ../JNW_TR_SKY130A
timestamp 1755333658
transform 1 0 3800 0 1 300
box 0 0 1880 3440
use JNWBIAS_OTACM  xad6
timestamp 1755440240
transform 1 0 8400 0 1 0
box 0 0 6800 10000
use JNWATR_PCH_4C5F0  xca1
timestamp 1740610800
transform 1 0 384 0 1 6100
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xca2
timestamp 1740610800
transform 1 0 384 0 1 6900
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xca3_0
timestamp 1740610800
transform 1 0 384 0 1 4500
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xca3_1
timestamp 1740610800
transform 1 0 384 0 1 5300
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xca3_2
timestamp 1740610800
transform 1 0 384 0 1 7700
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xca3_3
timestamp 1740610800
transform 1 0 384 0 1 8500
box -184 -128 1336 928
use JNWTR_CAPX1  xd1_0
timestamp 1737500400
transform 1 0 6500 0 1 5200
box 0 0 1080 1080
use JNWBIAS_BIPOLAR  xe1
timestamp 1755432682
transform 1 0 4217 0 1 4817
box -117 -117 4317 4317
use JNWTR_RPPO4  xf1
timestamp 1755333658
transform -1 0 3680 0 1 300
box 0 0 1880 3440
use JNWATR_NCH_4C5F0  xg7
timestamp 1740610800
transform 1 0 384 0 1 740
box -184 -128 1336 928
use JNWATR_NCH_4CTAPBOT  XJNWATR_NCH_4CTAPBOT2 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 384 0 1 260
box -184 -128 1336 608
use JNWATR_NCH_4CTAPTOP  XJNWATR_NCH_4CTAPTOP3 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 384 0 1 3140
box -184 -128 1336 608
use JNWATR_PCH_4CTAPBOT  XJNWATR_PCH_4CTAPBOT0
timestamp 1740610800
transform -1 0 1536 0 1 4039
box -184 -128 1336 608
use JNWATR_PCH_4CTAPTOP  XJNWATR_PCH_4CTAPTOP1
timestamp 1740610800
transform 1 0 384 0 1 9300
box -184 -128 1336 608
<< labels >>
flabel metal2 s 4095 6624 4287 6816 0 FreeSans 1600 0 0 0 VD1
flabel metal2 s 4231 7332 4423 7524 0 FreeSans 1600 0 0 0 VR1
flabel locali s 0 2 3046 400 0 FreeSans 1600 0 0 0 VSS
port 19 nsew
flabel locali s 0 9420 1632 10000 0 FreeSans 1600 0 0 0 VDD_1V8
port 17 nsew
flabel metal1 s 14352 9024 14544 9216 0 FreeSans 1600 0 0 0 LPI
port 16 nsew
flabel metal1 s 14352 8564 14544 8756 0 FreeSans 1600 0 0 0 LPO
port 15 nsew
flabel metal2 1664 3584 1856 3776 0 FreeSans 1600 0 0 0 VD2
flabel metal2 4564 3924 4756 4116 0 FreeSans 1600 0 0 0 VR1
flabel metal1 s 540 2000 604 2064 0 FreeSans 1600 0 0 0 STARTUP_1V8
port 14 nsew
flabel metal2 s 4 8676 1456 8868 0 FreeSans 1600 0 0 0 IBP_1U[1]
port 5 nsew
flabel metal2 s 4 7804 1456 7996 0 FreeSans 1600 0 0 0 IBP_1U[0]
port 6 nsew
flabel metal2 s 4 5404 1456 5596 0 FreeSans 1600 0 0 0 IBP_1U[2]
port 7 nsew
flabel metal2 s 4 4604 1456 4796 0 FreeSans 1600 0 0 0 IBP_1U[3]
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 15200 10000
<< end >>
