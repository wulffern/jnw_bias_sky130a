magic
tech sky130A
timestamp 1756046330
<< locali >>
rect 0 4935 3400 5000
rect 0 4915 1179 4935
rect 0 4825 347 4915
rect 437 4845 1179 4915
rect 1269 4927 3400 4935
rect 1269 4845 2193 4927
rect 437 4825 2193 4845
rect 0 4813 2193 4825
rect 2307 4813 3400 4927
rect 0 4800 3400 4813
rect 1000 4400 1100 4800
rect 290 4020 420 4060
rect 2350 2750 2450 2950
rect 2170 2020 2310 2060
rect 2740 2020 2880 2060
rect 2160 1620 2300 1660
rect 2730 1620 2870 1660
rect 2160 1220 2300 1260
rect 2730 1220 2870 1260
rect 2170 820 2310 860
rect 2740 820 2880 860
rect 2600 200 2700 500
rect 0 145 3400 200
rect 0 55 2211 145
rect 2301 55 2787 145
rect 2877 55 3400 145
rect 0 0 3400 55
<< viali >>
rect 347 4825 437 4915
rect 1179 4845 1269 4935
rect 2193 4813 2307 4927
rect 2190 4360 2310 4480
rect 2655 4375 2745 4465
rect 2211 55 2301 145
rect 2787 55 2877 145
<< metal1 >>
rect 1176 4935 1272 4941
rect 344 4915 440 4921
rect 344 4825 347 4915
rect 437 4825 440 4915
rect 281 4234 284 4266
rect 316 4234 319 4266
rect 284 4174 316 4234
rect 344 4072 440 4825
rect 1176 4845 1179 4935
rect 1269 4845 1272 4935
rect 1112 4266 1144 4269
rect 1112 4164 1144 4234
rect 1176 4042 1272 4845
rect 2190 4927 2310 4933
rect 2190 4813 2193 4927
rect 2307 4813 2310 4927
rect 2190 4490 2310 4813
rect 2180 4480 2330 4490
rect 2180 4360 2190 4480
rect 2310 4360 2330 4480
rect 2640 4465 2790 4500
rect 2640 4375 2655 4465
rect 2745 4375 2790 4465
rect 2640 4360 2790 4375
rect 2180 4350 2330 4360
rect 1622 4198 1718 4201
rect 1622 4099 1718 4102
rect 792 4008 888 4011
rect 792 3909 888 3912
rect 2400 4008 2496 4011
rect 342 3820 438 3823
rect 280 694 312 3756
rect 1170 3820 1290 3830
rect 438 3724 440 3818
rect 342 3721 440 3724
rect 344 3608 440 3721
rect 356 868 440 3544
rect 792 1830 888 3758
rect 1170 3724 1176 3820
rect 1272 3724 1290 3820
rect 1170 3720 1290 3724
rect 1176 3712 1256 3720
rect 1176 3572 1272 3712
rect 780 1818 900 1830
rect 780 1722 792 1818
rect 888 1722 900 1818
rect 780 1710 900 1722
rect 792 802 888 1710
rect 1112 684 1144 3546
rect 1178 936 1262 3572
rect 1624 1080 1720 3820
rect 2400 2456 2496 3912
rect 2652 3820 2748 4360
rect 2652 3721 2748 3724
rect 2976 4198 3072 4201
rect 1610 1068 1730 1080
rect 1610 972 1624 1068
rect 1720 972 1730 1068
rect 1610 960 1730 972
rect 1624 902 1720 960
rect 2144 634 2176 2366
rect 2208 145 2304 2448
rect 2400 1821 2496 2008
rect 2400 1818 2498 1821
rect 2400 1722 2402 1818
rect 2400 1719 2498 1722
rect 2400 862 2496 1719
rect 2720 934 2752 2396
rect 2208 55 2211 145
rect 2301 55 2304 145
rect 2208 49 2304 55
rect 2784 145 2880 2548
rect 2976 2522 3072 4102
rect 2976 1071 3072 2024
rect 2972 1068 3072 1071
rect 3068 972 3072 1068
rect 2972 969 3072 972
rect 2976 872 3072 969
rect 2784 55 2787 145
rect 2877 55 2880 145
rect 2784 49 2880 55
<< via1 >>
rect 284 4234 316 4266
rect 1112 4234 1144 4266
rect 1622 4102 1718 4198
rect 792 3912 888 4008
rect 2400 3912 2496 4008
rect 342 3724 438 3820
rect 1176 3724 1272 3820
rect 792 1722 888 1818
rect 2652 3724 2748 3820
rect 2976 4102 3072 4198
rect 1624 972 1720 1068
rect 2402 1722 2498 1818
rect 2972 972 3068 1068
<< metal2 >>
rect 284 4266 316 4269
rect 316 4234 1112 4266
rect 1144 4234 1147 4266
rect 284 4231 316 4234
rect 1619 4102 1622 4198
rect 1718 4102 2976 4198
rect 3072 4102 3075 4198
rect 789 3912 792 4008
rect 888 3912 2400 4008
rect 2496 3912 2499 4008
rect 1170 3820 1290 3830
rect 339 3724 342 3820
rect 438 3724 1176 3820
rect 1272 3724 2652 3820
rect 2748 3724 2751 3820
rect 1170 3720 1290 3724
rect 780 1818 900 1830
rect 780 1722 792 1818
rect 888 1722 2402 1818
rect 2498 1722 2501 1818
rect 780 1710 900 1722
rect 1610 1068 1730 1080
rect 1610 972 1624 1068
rect 1720 972 2972 1068
rect 3068 972 3071 1068
rect 1610 960 1730 972
use JNWATR_PCH_12C1F2  xba1_0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 200 0 1 640
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xba1_1
timestamp 1740610800
transform 1 0 200 0 1 1040
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xba1_2
timestamp 1740610800
transform 1 0 200 0 1 1440
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xba1_3
timestamp 1740610800
transform 1 0 200 0 1 1840
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xba1_4
timestamp 1740610800
transform 1 0 200 0 1 2240
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xba1_5
timestamp 1740610800
transform 1 0 200 0 1 2640
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xba1_6
timestamp 1740610800
transform 1 0 200 0 1 3040
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xba1_7
timestamp 1740610800
transform 1 0 200 0 1 3440
box -92 -64 924 464
use JNWATR_PCH_12C5F0  xba6 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 200 0 1 3840
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xbb2_0
timestamp 1740610800
transform 1 0 1032 0 1 640
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xbb2_1
timestamp 1740610800
transform 1 0 1032 0 1 1040
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xbb2_2
timestamp 1740610800
transform 1 0 1032 0 1 1440
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xbb2_3
timestamp 1740610800
transform 1 0 1032 0 1 1840
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xbb2_4
timestamp 1740610800
transform 1 0 1032 0 1 2240
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xbb2_5
timestamp 1740610800
transform 1 0 1032 0 1 2640
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xbb2_6
timestamp 1740610800
transform 1 0 1032 0 1 3040
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xbb2_7
timestamp 1740610800
transform 1 0 1032 0 1 3440
box -92 -64 924 464
use JNWATR_PCH_12C5F0  xbb3
timestamp 1740610800
transform 1 0 1032 0 1 3840
box -92 -64 924 464
use JNWATR_NCH_4C5F0  xca1_0 JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 2064 0 1 640
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xca1_1
timestamp 1740610800
transform 1 0 2064 0 1 1040
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xca1_2
timestamp 1740610800
transform 1 0 2064 0 1 1440
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xca1_3
timestamp 1740610800
transform 1 0 2064 0 1 1840
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xca3
timestamp 1740610800
transform 1 0 2064 0 1 2240
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xcb2_0
timestamp 1740610800
transform 1 0 2640 0 1 640
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xcb2_1
timestamp 1740610800
transform 1 0 2640 0 1 1040
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xcb2_2
timestamp 1740610800
transform 1 0 2640 0 1 1440
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xcb2_3
timestamp 1740610800
transform 1 0 2640 0 1 1840
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xcb4
timestamp 1740610800
transform 1 0 2640 0 1 2240
box -92 -64 668 464
use JNWTR_RPPO4  xd2 JNW_TR_SKY130A
timestamp 1755333658
transform 1 0 2000 0 1 2900
box 0 0 940 1720
use JNWATR_NCH_4CTAPBOT  XJNWATR_NCH_4CTAPBOT4 JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 2064 0 1 400
box -92 -64 668 304
use JNWATR_NCH_4CTAPBOT  XJNWATR_NCH_4CTAPBOT6
timestamp 1740610800
transform 1 0 2640 0 1 400
box -92 -64 668 304
use JNWATR_NCH_4CTAPTOP  XJNWATR_NCH_4CTAPTOP5 JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 2064 0 1 2640
box -92 -64 668 304
use JNWATR_NCH_4CTAPTOP  XJNWATR_NCH_4CTAPTOP7
timestamp 1740610800
transform 1 0 2640 0 1 2640
box -92 -64 668 304
use JNWATR_PCH_12CTAPBOT  XJNWATR_PCH_12CTAPBOT0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 200 0 1 400
box -92 -64 924 304
use JNWATR_PCH_12CTAPBOT  XJNWATR_PCH_12CTAPBOT2
timestamp 1740610800
transform 1 0 1032 0 1 400
box -92 -64 924 304
use JNWATR_PCH_12CTAPTOP  XJNWATR_PCH_12CTAPTOP1 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 200 0 1 4240
box -92 -64 924 304
use JNWATR_PCH_12CTAPTOP  XJNWATR_PCH_12CTAPTOP3
timestamp 1740610800
transform 1 0 1032 0 1 4240
box -92 -64 924 304
<< labels >>
flabel locali 0 4800 347 5000 0 FreeSans 800 0 0 0 VDD_1V8
port 0 nsew
flabel locali 0 0 2211 200 0 FreeSans 800 0 0 0 VSS
port 1 nsew
flabel metal1 280 694 312 3756 0 FreeSans 800 0 0 0 VIN
port 2 nsew
flabel metal1 1112 684 1144 3546 0 FreeSans 800 0 0 0 VIP
port 3 nsew
flabel metal1 2976 2522 3072 4102 0 FreeSans 800 0 0 0 VO
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 3400 5000
<< end >>
