magic
tech sky130A
magscale 1 2
timestamp 1756159200
<< checkpaint >>
rect 0 0 28854 10320
<< metal3 >>
rect 8652 4874 12452 5074
rect 9092 4434 9292 9594
rect 10452 4434 10652 9594
rect 11812 4434 12012 9594
rect 8652 6234 12452 6434
rect 9092 4434 9292 9594
rect 10452 4434 10652 9594
rect 11812 4434 12012 9594
rect 8652 7594 12452 7794
rect 9092 4434 9292 9594
rect 10452 4434 10652 9594
rect 11812 4434 12012 9594
rect 8652 8954 9732 9154
rect 9092 4434 9292 9594
<< metal4 >>
rect 8652 4874 12452 5074
rect 9092 4434 9292 9594
rect 10452 4434 10652 9594
rect 11812 4434 12012 9594
rect 8652 6234 12452 6434
rect 9092 4434 9292 9594
rect 10452 4434 10652 9594
rect 11812 4434 12012 9594
rect 8652 7594 12452 7794
rect 9092 4434 9292 9594
rect 10452 4434 10652 9594
rect 11812 4434 12012 9594
rect 8652 8954 9732 9154
rect 9092 4434 9292 9594
use JNWBIAS_OTACM xaota6 ../JNW_BIAS_SKY130A
transform 1 0 0 0 1 0
box 0 0 6800 10000
use JNWATR_PCH_4C5F0 xb1<0> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 0
box 7100 0 8252 800
use JNWATR_PCH_4C5F0 xb1<1> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 800
box 7100 800 8252 1600
use JNWATR_PCH_4C5F0 xb1<2> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 1600
box 7100 1600 8252 2400
use JNWATR_PCH_4C5F0 xb1<3> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 2400
box 7100 2400 8252 3200
use JNWATR_PCH_4C5F0 xb3<0> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 3200
box 7100 3200 8252 4000
use JNWATR_PCH_4C5F0 xb3<1> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 4000
box 7100 4000 8252 4800
use JNWATR_PCH_4C5F0 xb3<2> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 4800
box 7100 4800 8252 5600
use JNWATR_PCH_4C5F0 xb3<3> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 5600
box 7100 5600 8252 6400
use JNWATR_PCH_4C5F0 xb7<0> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 6400
box 7100 6400 8252 7200
use JNWATR_PCH_4C5F0 xb7<1> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 7200
box 7100 7200 8252 8000
use JNWATR_PCH_4C5F0 xb7<2> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 8000
box 7100 8000 8252 8800
use JNWATR_PCH_4C5F0 xb7<3> ../JNW_ATR_SKY130A
transform 1 0 7100 0 1 8800
box 7100 8800 8252 9600
use JNWBIAS_BIPOLAR xbc1 ../JNW_BIAS_SKY130A
transform 1 0 8652 0 1 0
box 8652 0 13086 4434
use JNWTR_CAPX1 xbc2<0> ../JNW_TR_SKY130A
transform 1 0 8652 0 1 4434
box 8652 4434 9732 5514
use JNWTR_CAPX1 xbc2<1> ../JNW_TR_SKY130A
transform 1 0 10012 0 1 4434
box 10012 4434 11092 5514
use JNWTR_CAPX1 xbc2<2> ../JNW_TR_SKY130A
transform 1 0 11372 0 1 4434
box 11372 4434 12452 5514
use JNWTR_CAPX1 xbc2<3> ../JNW_TR_SKY130A
transform 1 0 8652 0 1 5794
box 8652 5794 9732 6874
use JNWTR_CAPX1 xbc2<4> ../JNW_TR_SKY130A
transform 1 0 10012 0 1 5794
box 10012 5794 11092 6874
use JNWTR_CAPX1 xbc2<5> ../JNW_TR_SKY130A
transform 1 0 11372 0 1 5794
box 11372 5794 12452 6874
use JNWTR_CAPX1 xbc2<6> ../JNW_TR_SKY130A
transform 1 0 8652 0 1 7154
box 8652 7154 9732 8234
use JNWTR_CAPX1 xbc2<7> ../JNW_TR_SKY130A
transform 1 0 10012 0 1 7154
box 10012 7154 11092 8234
use JNWTR_CAPX1 xbc2<8> ../JNW_TR_SKY130A
transform 1 0 11372 0 1 7154
box 11372 7154 12452 8234
use JNWTR_CAPX1 xbc2<9> ../JNW_TR_SKY130A
transform 1 0 8652 0 1 8514
box 8652 8514 9732 9594
use JNWTR_RPPO8 xc11 ../JNW_TR_SKY130A
transform 1 0 13386 0 1 0
box 13386 0 16130 3440
use JNWTR_RPPO16 xc12 ../JNW_TR_SKY130A
transform 1 0 13386 0 1 3440
box 13386 3440 17858 6880
use JNWTR_RPPO16 xc9 ../JNW_TR_SKY130A
transform 1 0 13386 0 1 6880
box 13386 6880 17858 10320
use JNWTR_RPPO8 xd10 ../JNW_TR_SKY130A
transform 1 0 18158 0 1 0
box 18158 0 20902 3440
use JNWTR_RPPO16 xd13 ../JNW_TR_SKY130A
transform 1 0 18158 0 1 3440
box 18158 3440 22630 6880
use JNWTR_RPPO16 xd7 ../JNW_TR_SKY130A
transform 1 0 18158 0 1 6880
box 18158 6880 22630 10320
use JNWTR_RPPO4 xe2 ../JNW_TR_SKY130A
transform 1 0 22930 0 1 0
box 22930 0 24810 3440
use JNWTR_RPPO16 xe3 ../JNW_TR_SKY130A
transform 1 0 22930 0 1 3440
box 22930 3440 27402 6880
use JNWTR_RPPO2 xe8 ../JNW_TR_SKY130A
transform 1 0 22930 0 1 6880
box 22930 6880 24378 10320
use JNWATR_NCH_4C5F0 xf4 ../JNW_ATR_SKY130A
transform 1 0 27702 0 1 0
box 27702 0 28854 800
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 28854 10320
<< end >>
