magic
tech sky130A
magscale 1 2
timestamp 1755336416
<< locali >>
rect -800 10200 10000 10600
rect -800 -200 -400 10200
rect 3600 8400 4000 10200
rect 6800 9600 7200 10200
rect 9600 7600 10000 10200
rect 8000 7200 10000 7600
rect -200 3600 9400 4000
rect 600 -200 1000 100
rect 2200 -200 2600 100
rect 9600 -200 10000 7200
rect -800 -600 10000 -200
use JNWTR_RPPO4  xab3 ../JNW_TR_SKY130A
timestamp 1755333658
transform 1 0 -200 0 1 0
box 0 0 1880 3440
use JNWTR_RPPO2  xac2 ../JNW_TR_SKY130A
timestamp 1755255778
transform 1 0 1800 0 1 0
box 0 0 1448 3440
use JNWBIAS_OTAR  xad6
timestamp 1755336416
transform 1 0 3500 0 1 0
box -100 -400 5800 3800
use JNWATR_PCH_4C5F0  xca1 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 -16 0 1 4808
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xca2
timestamp 1740610800
transform 1 0 -16 0 1 5608
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xca3_0
timestamp 1740610800
transform 1 0 -16 0 1 6408
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xca3_1
timestamp 1740610800
transform 1 0 -16 0 1 7208
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xca3_2
timestamp 1740610800
transform 1 0 -16 0 1 8008
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xca3_3
timestamp 1740610800
transform 1 0 -16 0 1 8808
box -184 -128 1336 928
use JNWTR_CAPX1  xd1_0 ../JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 8184 0 1 4208
box 0 0 1080 1080
use JNWTR_CAPX1  xd1_1
timestamp 1737500400
transform 1 0 8184 0 1 5688
box 0 0 1080 1080
use JNWBIAS_BIPOLAR  xe1
timestamp 1755335025
transform 1 0 1701 0 1 4405
box -117 -117 4317 4317
use JNWTR_RPPO4  xf1
timestamp 1755333658
transform 1 0 6184 0 1 4288
box 0 0 1880 3440
use JNWATR_NCH_4C5F0  xg7 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 6368 0 1 8616
box -184 -128 1336 928
use JNWATR_NCH_4CTAPBOT  XJNWATR_NCH_4CTAPBOT2 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 6368 0 1 8136
box -184 -128 1336 608
use JNWATR_NCH_4CTAPTOP  XJNWATR_NCH_4CTAPTOP3 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 6368 0 1 9416
box -184 -128 1336 608
use JNWATR_PCH_4CTAPBOT  XJNWATR_PCH_4CTAPBOT0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 -16 0 1 4328
box -184 -128 1336 608
use JNWATR_PCH_4CTAPTOP  XJNWATR_PCH_4CTAPTOP1 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 -16 0 1 9608
box -184 -128 1336 608
<< properties >>
string FIXED_BBOX 0 0 10818 9800
<< end >>
