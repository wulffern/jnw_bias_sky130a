magic
tech sky130A
timestamp 1755432610
<< locali >>
rect -200 4535 3200 4600
rect -200 4515 979 4535
rect -200 4425 147 4515
rect 237 4445 979 4515
rect 1069 4527 3200 4535
rect 1069 4445 1993 4527
rect 237 4425 1993 4445
rect -200 4413 1993 4425
rect 2107 4413 3200 4527
rect -200 4400 3200 4413
rect 800 4000 900 4400
rect 90 3620 220 3660
rect 2150 2350 2250 2550
rect 1970 1620 2110 1660
rect 2540 1620 2680 1660
rect 1960 1220 2100 1260
rect 2530 1220 2670 1260
rect 1960 820 2100 860
rect 2530 820 2670 860
rect 1970 420 2110 460
rect 2540 420 2680 460
rect 2400 -200 2500 100
rect -200 -255 3200 -200
rect -200 -345 2011 -255
rect 2101 -345 2587 -255
rect 2677 -345 3200 -255
rect -200 -400 3200 -345
<< viali >>
rect 147 4425 237 4515
rect 979 4445 1069 4535
rect 1993 4413 2107 4527
rect 1990 3960 2110 4080
rect 2455 3975 2545 4065
rect 2011 -345 2101 -255
rect 2587 -345 2677 -255
<< metal1 >>
rect 976 4535 1072 4541
rect 144 4515 240 4521
rect 144 4425 147 4515
rect 237 4425 240 4515
rect 81 3834 84 3866
rect 116 3834 119 3866
rect 84 3774 116 3834
rect 144 3672 240 4425
rect 976 4445 979 4535
rect 1069 4445 1072 4535
rect 912 3866 944 3869
rect 912 3764 944 3834
rect 976 3642 1072 4445
rect 1990 4527 2110 4533
rect 1990 4413 1993 4527
rect 2107 4413 2110 4527
rect 1990 4090 2110 4413
rect 1980 4080 2130 4090
rect 1980 3960 1990 4080
rect 2110 3960 2130 4080
rect 2440 4065 2590 4100
rect 2440 3975 2455 4065
rect 2545 3975 2590 4065
rect 2440 3960 2590 3975
rect 1980 3950 2130 3960
rect 1422 3798 1518 3801
rect 1422 3699 1518 3702
rect 592 3608 688 3611
rect 592 3509 688 3512
rect 2200 3608 2296 3611
rect 142 3420 238 3423
rect 80 294 112 3356
rect 970 3420 1090 3430
rect 238 3324 240 3418
rect 142 3321 240 3324
rect 144 3208 240 3321
rect 156 468 240 3144
rect 592 1430 688 3358
rect 970 3324 976 3420
rect 1072 3324 1090 3420
rect 970 3320 1090 3324
rect 976 3312 1056 3320
rect 976 3172 1072 3312
rect 580 1418 700 1430
rect 580 1322 592 1418
rect 688 1322 700 1418
rect 580 1310 700 1322
rect 592 402 688 1310
rect 912 284 944 3146
rect 978 536 1062 3172
rect 1424 680 1520 3420
rect 2200 2056 2296 3512
rect 2452 3420 2548 3960
rect 2452 3321 2548 3324
rect 2776 3798 2872 3801
rect 1410 668 1530 680
rect 1410 572 1424 668
rect 1520 572 1530 668
rect 1410 560 1530 572
rect 1424 502 1520 560
rect 1944 234 1976 1966
rect 2008 -255 2104 2048
rect 2200 1421 2296 1608
rect 2200 1418 2298 1421
rect 2200 1322 2202 1418
rect 2200 1319 2298 1322
rect 2200 462 2296 1319
rect 2520 534 2552 1996
rect 2008 -345 2011 -255
rect 2101 -345 2104 -255
rect 2008 -351 2104 -345
rect 2584 -255 2680 2148
rect 2776 2122 2872 3702
rect 2776 671 2872 1624
rect 2772 668 2872 671
rect 2868 572 2872 668
rect 2772 569 2872 572
rect 2776 472 2872 569
rect 2584 -345 2587 -255
rect 2677 -345 2680 -255
rect 2584 -351 2680 -345
<< via1 >>
rect 84 3834 116 3866
rect 912 3834 944 3866
rect 1422 3702 1518 3798
rect 592 3512 688 3608
rect 2200 3512 2296 3608
rect 142 3324 238 3420
rect 976 3324 1072 3420
rect 592 1322 688 1418
rect 2452 3324 2548 3420
rect 2776 3702 2872 3798
rect 1424 572 1520 668
rect 2202 1322 2298 1418
rect 2772 572 2868 668
<< metal2 >>
rect 84 3866 116 3869
rect 116 3834 912 3866
rect 944 3834 947 3866
rect 84 3831 116 3834
rect 1419 3702 1422 3798
rect 1518 3702 2776 3798
rect 2872 3702 2875 3798
rect 589 3512 592 3608
rect 688 3512 2200 3608
rect 2296 3512 2299 3608
rect 970 3420 1090 3430
rect 139 3324 142 3420
rect 238 3324 976 3420
rect 1072 3324 2452 3420
rect 2548 3324 2551 3420
rect 970 3320 1090 3324
rect 580 1418 700 1430
rect 580 1322 592 1418
rect 688 1322 2202 1418
rect 2298 1322 2301 1418
rect 580 1310 700 1322
rect 1410 668 1530 680
rect 1410 572 1424 668
rect 1520 572 2772 668
rect 2868 572 2871 668
rect 1410 560 1530 572
use JNWATR_PCH_12C1F2  xba1_0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 0 0 1 240
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xba1_1
timestamp 1740610800
transform 1 0 0 0 1 640
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xba1_2
timestamp 1740610800
transform 1 0 0 0 1 1040
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xba1_3
timestamp 1740610800
transform 1 0 0 0 1 1440
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xba1_4
timestamp 1740610800
transform 1 0 0 0 1 1840
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xba1_5
timestamp 1740610800
transform 1 0 0 0 1 2240
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xba1_6
timestamp 1740610800
transform 1 0 0 0 1 2640
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xba1_7
timestamp 1740610800
transform 1 0 0 0 1 3040
box -92 -64 924 464
use JNWATR_PCH_12C5F0  xba6 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 0 0 1 3440
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xbb2_0
timestamp 1740610800
transform 1 0 832 0 1 240
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xbb2_1
timestamp 1740610800
transform 1 0 832 0 1 640
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xbb2_2
timestamp 1740610800
transform 1 0 832 0 1 1040
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xbb2_3
timestamp 1740610800
transform 1 0 832 0 1 1440
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xbb2_4
timestamp 1740610800
transform 1 0 832 0 1 1840
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xbb2_5
timestamp 1740610800
transform 1 0 832 0 1 2240
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xbb2_6
timestamp 1740610800
transform 1 0 832 0 1 2640
box -92 -64 924 464
use JNWATR_PCH_12C1F2  xbb2_7
timestamp 1740610800
transform 1 0 832 0 1 3040
box -92 -64 924 464
use JNWATR_PCH_12C5F0  xbb3
timestamp 1740610800
transform 1 0 832 0 1 3440
box -92 -64 924 464
use JNWATR_NCH_4C5F0  xca1_0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 1864 0 1 240
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xca1_1
timestamp 1740610800
transform 1 0 1864 0 1 640
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xca1_2
timestamp 1740610800
transform 1 0 1864 0 1 1040
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xca1_3
timestamp 1740610800
transform 1 0 1864 0 1 1440
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xca3
timestamp 1740610800
transform 1 0 1864 0 1 1840
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xcb2_0
timestamp 1740610800
transform 1 0 2440 0 1 240
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xcb2_1
timestamp 1740610800
transform 1 0 2440 0 1 640
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xcb2_2
timestamp 1740610800
transform 1 0 2440 0 1 1040
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xcb2_3
timestamp 1740610800
transform 1 0 2440 0 1 1440
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xcb4
timestamp 1740610800
transform 1 0 2440 0 1 1840
box -92 -64 668 464
use JNWTR_RPPO4  xd2 ../JNW_TR_SKY130A
timestamp 1755333658
transform 1 0 1800 0 1 2500
box 0 0 940 1720
use JNWATR_NCH_4CTAPBOT  XJNWATR_NCH_4CTAPBOT4 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 1864 0 1 0
box -92 -64 668 304
use JNWATR_NCH_4CTAPBOT  XJNWATR_NCH_4CTAPBOT6
timestamp 1740610800
transform 1 0 2440 0 1 0
box -92 -64 668 304
use JNWATR_NCH_4CTAPTOP  XJNWATR_NCH_4CTAPTOP5 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 1864 0 1 2240
box -92 -64 668 304
use JNWATR_NCH_4CTAPTOP  XJNWATR_NCH_4CTAPTOP7
timestamp 1740610800
transform 1 0 2440 0 1 2240
box -92 -64 668 304
use JNWATR_PCH_12CTAPBOT  XJNWATR_PCH_12CTAPBOT0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 0 0 1 0
box -92 -64 924 304
use JNWATR_PCH_12CTAPBOT  XJNWATR_PCH_12CTAPBOT2
timestamp 1740610800
transform 1 0 832 0 1 0
box -92 -64 924 304
use JNWATR_PCH_12CTAPTOP  XJNWATR_PCH_12CTAPTOP1 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 0 0 1 3840
box -92 -64 924 304
use JNWATR_PCH_12CTAPTOP  XJNWATR_PCH_12CTAPTOP3
timestamp 1740610800
transform 1 0 832 0 1 3840
box -92 -64 924 304
<< labels >>
flabel locali -200 4400 147 4600 0 FreeSans 800 0 0 0 VDD_1V8
port 0 nsew
flabel locali -200 -400 2011 -200 0 FreeSans 800 0 0 0 VSS
port 1 nsew
flabel metal1 80 294 112 3356 0 FreeSans 800 0 0 0 VIN
port 2 nsew
flabel metal1 912 284 944 3146 0 FreeSans 800 0 0 0 VIP
port 3 nsew
flabel metal1 2776 2056 2872 3702 0 FreeSans 800 0 0 0 VO
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 4156 4080
<< end >>
