magic
tech sky130A
magscale 1 2
timestamp 1755339872
<< locali >>
rect -800 10200 10000 10600
rect -800 -200 -400 10200
rect 3600 8400 4000 10200
rect 6800 9600 7200 10200
rect 9600 7600 10000 10200
rect 8000 7448 10000 7600
rect 6504 7390 6848 7396
rect 6504 7210 6662 7390
rect 6842 7210 6848 7390
rect 6504 7204 6848 7210
rect 7460 7208 10000 7448
rect 8000 7200 10000 7208
rect 300 4000 700 4600
rect -200 3969 9400 4000
rect -200 3910 7271 3969
rect -200 3730 730 3910
rect 910 3730 7271 3910
rect -200 3600 7271 3730
rect 6765 3591 7271 3600
rect 7649 3600 9400 3969
rect 7649 3591 7655 3600
rect 6765 3585 7655 3591
rect 600 -200 1000 100
rect 2200 -200 2600 100
rect 9600 -200 10000 7200
rect -800 -212 10000 -200
rect -800 -600 2240 -212
rect 2640 -600 10000 -212
<< viali >>
rect 6662 7210 6842 7390
rect 730 3730 910 3910
rect 7271 3591 7649 3969
rect 230 2970 410 3150
rect 1088 2920 1316 3160
rect 2106 2926 2334 3154
rect 2600 2920 2840 3160
rect 2240 -600 2640 -212
<< metal1 >>
rect 138 9768 144 9832
rect 208 9768 214 9832
rect 144 5428 208 9768
rect 272 7036 464 9196
rect 650 8984 656 9176
rect 848 8984 854 9176
rect 6528 8708 6592 10592
rect 8955 9885 9325 9891
rect 7168 9832 7232 9838
rect 7168 9268 7232 9768
rect 650 8104 656 8296
rect 848 8104 854 8296
rect 640 7832 860 7840
rect 640 7640 656 7832
rect 848 7640 860 7832
rect 640 7620 860 7640
rect 1240 7832 1480 7860
rect 1240 7640 1264 7832
rect 1456 7640 1480 7832
rect 1240 7620 1480 7640
rect 272 4924 464 6844
rect 464 3916 656 3922
rect 656 3910 922 3916
rect 656 3730 730 3910
rect 910 3730 922 3910
rect 656 3724 922 3730
rect 464 3718 656 3724
rect 224 3536 416 3542
rect 224 3150 416 3344
rect 1264 3536 1456 7620
rect 6656 7390 6848 8996
rect 6656 7210 6662 7390
rect 6842 7210 6848 7390
rect 6656 7198 6848 7210
rect 3604 6776 3796 6782
rect 3604 6578 3796 6584
rect 1264 3338 1456 3344
rect 2600 3180 2840 4880
rect 7665 3975 8055 3981
rect 7259 3969 7665 3975
rect 7259 3591 7271 3969
rect 7649 3591 7665 3969
rect 7259 3585 7665 3591
rect 7665 3579 8055 3585
rect 224 2970 230 3150
rect 410 2970 416 3150
rect 224 2036 416 2970
rect 1082 3160 1322 3172
rect 2580 3160 2860 3180
rect 1082 2920 1088 3160
rect 1316 3154 2346 3160
rect 1316 2926 2106 3154
rect 2334 2926 2346 3154
rect 1316 2920 2346 2926
rect 2580 2920 2600 3160
rect 2840 2920 2860 3160
rect 1082 2908 1322 2920
rect 2580 2900 2860 2920
rect 8955 2845 9325 9515
rect 224 1844 5756 2036
rect 2240 1520 2640 1526
rect 2240 -206 2640 1120
rect 5364 1136 5556 1142
rect 5556 944 5736 1136
rect 8955 955 9325 2475
rect 5364 938 5556 944
rect 2228 -212 2652 -206
rect 2228 -600 2240 -212
rect 2640 -600 2652 -212
rect 2228 -606 2652 -600
<< via1 >>
rect 144 9768 208 9832
rect 656 8984 848 9176
rect 7168 9768 7232 9832
rect 8955 9515 9325 9885
rect 656 8104 848 8296
rect 656 7640 848 7832
rect 1264 7640 1456 7832
rect 272 6844 464 7036
rect 656 6584 848 6776
rect 656 5704 848 5896
rect 656 4904 848 5096
rect 464 3724 656 3916
rect 224 3344 416 3536
rect 3604 6584 3796 6776
rect 1264 3344 1456 3536
rect 7665 3585 8055 3975
rect 2240 1120 2640 1520
rect 5364 944 5556 1136
<< metal2 >>
rect 55 9900 8909 9905
rect 55 9832 8544 9900
rect 55 9768 144 9832
rect 208 9768 7168 9832
rect 7232 9768 8544 9832
rect 55 9540 8544 9768
rect 8904 9885 8913 9900
rect 8904 9540 8955 9885
rect 55 9535 8955 9540
rect 8015 9515 8955 9535
rect 9325 9515 9331 9885
rect 656 9176 848 9182
rect -796 8984 656 9176
rect 656 8978 848 8984
rect 656 8300 848 8302
rect 640 8296 860 8300
rect -796 8104 656 8296
rect 848 8104 860 8296
rect 640 8080 860 8104
rect 640 7832 860 7840
rect 1240 7832 1480 7860
rect 640 7640 656 7832
rect 848 7640 1264 7832
rect 1456 7640 1480 7832
rect 640 7620 860 7640
rect 1240 7620 1480 7640
rect 260 7036 480 7040
rect 260 6844 272 7036
rect 464 6844 480 7036
rect 260 6840 480 6844
rect 272 6766 464 6840
rect 272 6575 464 6584
rect 640 6776 860 6780
rect 640 6584 656 6776
rect 848 6584 3104 6776
rect 3296 6584 3604 6776
rect 3796 6584 3802 6776
rect 640 6560 860 6584
rect 660 5896 880 5920
rect -796 5704 656 5896
rect 848 5704 880 5896
rect 660 5700 880 5704
rect 640 5096 860 5100
rect -796 4904 656 5096
rect 848 4904 860 5096
rect 640 4880 860 4904
rect -800 3975 10000 4000
rect -800 3916 7665 3975
rect -800 3911 464 3916
rect -800 3729 277 3911
rect 459 3729 464 3911
rect -800 3724 464 3729
rect 656 3724 7665 3916
rect -800 3600 7665 3724
rect 7659 3585 7665 3600
rect 8055 3970 10000 3975
rect 8055 3590 8150 3970
rect 8530 3600 10000 3970
rect 8530 3590 8535 3600
rect 8055 3585 8535 3590
rect 8150 3581 8530 3585
rect 218 3344 224 3536
rect 416 3344 1264 3536
rect 1456 3344 1462 3536
rect 2139 1539 4001 2141
rect 2140 1520 2720 1539
rect 2140 1120 2240 1520
rect 2640 1120 2720 1520
rect 3104 1131 5364 1136
rect 2140 1100 2720 1120
rect 3100 949 3109 1131
rect 3291 949 5364 1131
rect 3104 944 5364 949
rect 5556 944 5562 1136
<< via2 >>
rect 8544 9540 8904 9900
rect 272 6584 464 6766
rect 3104 6584 3296 6776
rect 277 3729 459 3911
rect 8150 3590 8530 3970
rect 3109 949 3291 1131
<< metal3 >>
rect 8539 9900 8909 9905
rect 8539 9540 8544 9900
rect 8904 9540 8909 9900
rect 3099 6776 3301 6781
rect 267 6766 469 6771
rect 267 6584 272 6766
rect 464 6584 469 6766
rect 267 6579 469 6584
rect 3099 6584 3104 6776
rect 3296 6584 3301 6776
rect 3099 6579 3301 6584
rect 272 3911 464 6579
rect 272 3729 277 3911
rect 459 3729 464 3911
rect 272 3724 464 3729
rect 3104 1131 3296 6579
rect 8539 4563 8909 9540
rect 8145 3974 8915 3975
rect 8145 3970 8526 3974
rect 8145 3590 8150 3970
rect 8145 3586 8526 3590
rect 8914 3586 8920 3974
rect 8145 3585 8915 3586
rect 3104 949 3109 1131
rect 3291 949 3296 1131
rect 3104 944 3296 949
<< via3 >>
rect 8526 3970 8914 3974
rect 8526 3590 8530 3970
rect 8530 3590 8914 3970
rect 8526 3586 8914 3590
<< metal4 >>
rect 8525 3974 8915 9295
rect 8525 3586 8526 3974
rect 8914 3586 8915 3974
rect 8525 3585 8915 3586
use JNWTR_CAPX1 JNWTR_CAPX1_0 ../JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 8200 0 1 7000
box 0 0 1080 1080
use JNWTR_RPPO4 xab3 ../JNW_TR_SKY130A
timestamp 1755333658
transform -1 0 1680 0 1 0
box 0 0 1880 3440
use JNWTR_RPPO2 xac2 ../JNW_TR_SKY130A
timestamp 1755255778
transform -1 0 3248 0 1 0
box 0 0 1448 3440
use JNWBIAS_OTAR xad6 ../JNW_BIAS_SKY130A
timestamp 1755336416
transform 1 0 3500 0 1 0
box -100 -400 5800 3800
use JNWATR_PCH_4C5F0 xca1 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 -16 0 1 6408
box -184 -128 1336 928
use JNWATR_PCH_4C5F0 xca2 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 -16 0 1 7208
box -184 -128 1336 928
use JNWATR_PCH_4C5F0 xca3_0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 -16 0 1 4808
box -184 -128 1336 928
use JNWATR_PCH_4C5F0 xca3_1 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 -16 0 1 5608
box -184 -128 1336 928
use JNWATR_PCH_4C5F0 xca3_2 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 -16 0 1 8008
box -184 -128 1336 928
use JNWATR_PCH_4C5F0 xca3_3 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 -16 0 1 8808
box -184 -128 1336 928
use JNWTR_CAPX1 xd1_0 ../JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 8184 0 1 4208
box 0 0 1080 1080
use JNWTR_CAPX1 xd1_1 ../JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 8200 0 1 5600
box 0 0 1080 1080
use JNWBIAS_BIPOLAR xe1 ../JNW_BIAS_SKY130A
timestamp 1755335025
transform 1 0 1701 0 1 4405
box -117 -117 4317 4317
use JNWTR_RPPO4 xf1 ../JNW_TR_SKY130A
timestamp 1755333658
transform -1 0 8064 0 1 4288
box 0 0 1880 3440
use JNWATR_NCH_4C5F0 xg7 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 6368 0 1 8616
box -184 -128 1336 928
use JNWATR_NCH_4CTAPBOT XJNWATR_NCH_4CTAPBOT2 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 6368 0 1 8136
box -184 -128 1336 608
use JNWATR_NCH_4CTAPTOP XJNWATR_NCH_4CTAPTOP3 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 6368 0 1 9416
box -184 -128 1336 608
use JNWATR_PCH_4CTAPBOT XJNWATR_PCH_4CTAPBOT0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 -16 0 1 4328
box -184 -128 1336 608
use JNWATR_PCH_4CTAPTOP XJNWATR_PCH_4CTAPTOP1 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 -16 0 1 9608
box -184 -128 1336 608
<< labels >>
flabel metal2 s -796 8984 656 9176 0 FreeSans 1600 0 0 0 IBP_1U[0]
port 5 nsew
flabel metal2 s -796 8104 656 8296 0 FreeSans 1600 0 0 0 IBP_1U[1]
port 6 nsew
flabel metal2 s -796 5704 656 5896 0 FreeSans 1600 0 0 0 IBP_1U[2]
port 7 nsew
flabel metal2 s -796 4904 656 5096 0 FreeSans 1600 0 0 0 IBP_1U[3]
port 8 nsew
flabel metal1 s 8955 2845 9325 3215 0 FreeSans 1600 0 0 0 LPI
port 9 nsew
flabel metal1 s 8955 2095 9325 2465 0 FreeSans 1600 0 0 0 LPO
port 10 nsew
flabel metal2 s -600 3600 277 4000 0 FreeSans 1600 0 0 0 VDD_1V8
port 12 nsew
flabel locali s -800 -600 2240 -200 0 FreeSans 1600 0 0 0 VSS
port 13 nsew
flabel metal1 s 6528 10528 6592 10592 0 FreeSans 1600 0 0 0 STARTUP_1V8
port 14 nsew
flabel metal1 s 224 1844 416 2970 0 FreeSans 1600 0 0 0 VR1
flabel metal2 s 3291 944 5364 1136 0 FreeSans 1600 0 0 0 VD1
flabel metal1 s 2600 3160 2840 5405 0 FreeSans 1600 0 0 0 VD2
<< properties >>
string FIXED_BBOX 0 0 10818 9800
<< end >>
