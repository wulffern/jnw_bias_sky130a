magic
tech sky130A
timestamp 1755256143
<< locali >>
rect -50 1865 2900 1900
rect -50 1835 293 1865
rect 323 1835 2900 1865
rect -50 1800 2900 1835
rect 290 1382 326 1488
rect 1350 1150 1450 1800
rect 2260 820 2400 860
rect 2300 145 2420 150
rect 2300 55 2303 145
rect 2393 100 2420 145
rect 2393 55 2500 100
rect 2300 50 2500 55
rect 300 -100 400 50
rect 2400 -100 2500 50
rect -50 -200 2900 -100
<< viali >>
rect 293 1835 323 1865
rect 290 1488 326 1518
rect 365 1475 455 1565
rect 2303 55 2393 145
<< metal1 >>
rect 290 1865 326 1871
rect 290 1835 293 1865
rect 323 1835 326 1865
rect 290 1521 326 1835
rect 422 1568 518 1571
rect 359 1565 422 1568
rect 284 1518 332 1521
rect 284 1488 290 1518
rect 326 1488 332 1518
rect 284 1485 332 1488
rect 359 1475 365 1565
rect 359 1472 422 1475
rect 422 1469 518 1472
rect 1168 1568 1264 1571
rect 1100 890 1140 1020
rect 1168 822 1264 1472
rect 1610 1020 1720 1030
rect 1610 924 1616 1020
rect 1712 924 1720 1020
rect 1610 920 1720 924
rect 2500 1020 2610 1030
rect 2500 924 2502 1020
rect 2598 924 2610 1020
rect 2500 920 2610 924
rect 1100 490 1140 620
rect 1168 452 1264 818
rect 2236 534 2268 766
rect 1610 356 1720 360
rect 1610 260 1616 356
rect 1712 260 1720 356
rect 1610 250 1720 260
rect 2300 145 2396 798
rect 2492 472 2778 568
rect 2500 356 2610 360
rect 2500 260 2502 356
rect 2598 260 2610 356
rect 2500 250 2610 260
rect 2300 55 2303 145
rect 2393 55 2396 145
rect 2300 49 2396 55
<< via1 >>
rect 422 1565 518 1568
rect 422 1475 455 1565
rect 455 1475 518 1565
rect 422 1472 518 1475
rect 1168 1472 1264 1568
rect 1616 924 1712 1020
rect 2502 924 2598 1020
rect 1616 260 1712 356
rect 2502 260 2598 356
<< metal2 >>
rect 419 1472 422 1568
rect 518 1472 1168 1568
rect 1264 1472 1267 1568
rect 1610 1020 1720 1030
rect 2500 1020 2610 1030
rect 1610 924 1616 1020
rect 1712 924 2502 1020
rect 2598 924 2610 1020
rect 1610 920 1720 924
rect 2500 920 2610 924
rect 1610 356 1720 360
rect 2500 356 2610 360
rect 1610 260 1616 356
rect 1712 260 2502 356
rect 2598 260 2610 356
rect 1610 250 1720 260
rect 2500 250 2610 260
use JNWTR_RPPO2  xa1 ../JNW_TR_SKY130A
timestamp 1755255778
transform 1 0 0 0 1 0
box 0 0 724 1720
use JNWATR_PCH_12C5F0  xb1 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 1024 0 1 240
box -92 -64 924 464
use JNWATR_PCH_12C5F0  xb2
timestamp 1740610800
transform 1 0 1024 0 1 640
box -92 -64 924 464
use JNWATR_NCH_4C5F0  xc1 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 2156 0 1 240
box -92 -64 668 464
use JNWATR_NCH_4C5F0  xc2
timestamp 1740610800
transform 1 0 2156 0 1 640
box -92 -64 668 464
use JNWATR_NCH_4CTAPBOT  XJNWATR_NCH_4CTAPBOT2 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 2156 0 1 0
box -92 -64 668 304
use JNWATR_NCH_4CTAPTOP  XJNWATR_NCH_4CTAPTOP3 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 2156 0 1 1040
box -92 -64 668 304
use JNWATR_PCH_12CTAPBOT  XJNWATR_PCH_12CTAPBOT0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 1024 0 1 0
box -92 -64 924 304
use JNWATR_PCH_12CTAPTOP  XJNWATR_PCH_12CTAPTOP1 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 1024 0 1 1040
box -92 -64 924 304
<< labels >>
flabel locali -50 1800 2900 1900 0 FreeSans 800 0 0 0 VDD_1V8
port 0 nsew
flabel locali -50 -200 2900 -100 0 FreeSans 800 0 0 0 VSS
port 1 nsew
flabel metal1 2492 472 2778 568 0 FreeSans 800 0 0 0 VO
port 2 nsew
flabel metal1 1104 890 1136 1020 0 FreeSans 800 0 0 0 VIP
port 3 nsew
flabel metal1 1104 490 1136 620 0 FreeSans 800 0 0 0 VIN
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2732 1720
<< end >>
